//===============================================================================================================
// Module: tb.sv
// Author: Viacheslav Tarasov
// email: sl-engineer@protonmail.com
//===============================================================================================================

import cross_bar_pkg::*;

module tb();

// generate variable
genvar i;

//---------------------------------------------------------------------------------------------------------------
// clock
//---------------------------------------------------------------------------------------------------------------
logic   device_clk;                                               // device clock
initial device_clk = 1'b0;
always #2.5ns device_clk = ~device_clk;                           // 200 MHz

//---------------------------------------------------------------------------------------------------------------
// reset  
//---------------------------------------------------------------------------------------------------------------
bit resetn = 1'b1;

initial begin
    resetn = 1'b0;
    repeat (20) @(posedge device_clk);
    resetn = 1'b1;
end

//---------------------------------------------------------------------------------------------------------------
// signals  
//---------------------------------------------------------------------------------------------------------------
logic [MASTER_N - 1: 0] req;
logic [MASTER_N - 1: 0] grant;

//---------------------------------------------------------------------------------------------------------------
// DUT 
//---------------------------------------------------------------------------------------------------------------
cross_bar_rr_arbiter dut (
                          // clk and asynchronus negative reset
                          .clk     (device_clk),
                          .aresetn (resetn),

                          // req and grant interface
                          .req     (req),
                          .grant   (grant)
                         );

//---------------------------------------------------------------------------------------------------------------
// testbench body 
//---------------------------------------------------------------------------------------------------------------
initial begin: main
  req = {MASTER_N{1'b0}};
  
  wait (resetn);
  repeat (3) @(posedge device_clk);
  
  @(posedge device_clk);
  req[0] = 1;
  @(posedge device_clk);
  req[0] = 0;
  @(posedge device_clk);
  req[0] = 1;
  req[1] = 1;
  @(posedge device_clk);
  req[2] = 1;
  req[1] = 0;
  @(posedge device_clk);
  req[3] = 1;
  req[2] = 0;
  @(posedge device_clk);
  req[3] = 0;
  @(posedge device_clk);
  req[0] = 0;
  
  
  #1us;
  $display("\n\n\n\n");
  $display("Test passed!");
  $display("\n\n\n\n");
  $stop;
end  

initial #10 $display("\n\n\n\n");

endmodule

